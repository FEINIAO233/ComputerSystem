module and2x(input a,b,output r);
	assign r=a & b;
endmodule
